//  head info

module module_name(
    //  IO PORT DECLARATIONS

);

//=======================
//  PARAMETER DEFINITIONS
//=======================



//======================
//  VARIABLE DEFINITIONS
//======================



//===============
//  DESIGN CODING
//===============



endmodule
